interface mux_interface;
  
  logic clk;
  logic rst;
  logic [15:0][32:0] i;
  logic [3:0] s;
  logic [32:0] y;

endinterface
